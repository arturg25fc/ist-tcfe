.OP
R1 0 2 1001.783861
R2 3 2 2073.072177
R3 2 5 3117.913022
R4 5 0 4111.352423
R5 5 6 3104.598426
R6 4 7 2071.733607
R7 7 8 1043.430656
Vx 6 8 8.535665
Vfalsa 0 4 0.0
Hd 5 8 Vfalsa 8295.559623
Gb 6 3 2 5 0.007270
.END
